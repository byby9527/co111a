`ifndef or_nt
  `include "or_nt.v"
`endif
`define and_nt 1

module and_nt(input a, input b, output out);

    // Put your code here

endmodule 
