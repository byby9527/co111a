`ifndef dmux4way
  `include "dmux4way.v"
`endif
`define dmux8way 1

module dmux8way(
    input       in,
    input [2:0] select,
    output      a,
    output      b,
    output      c,
    output      d,
    output      e,
    output      f,
    output      g,
    output      h
);

    // Put your code here

endmodule
