`ifndef dmux
  `include "dmux.v"
`endif
`define dmux4way 1

module dmux4way(
    input       in,
    input [1:0] sel,
    output      a,
    output      b,
    output      c,
    output      d
);

    // Put your code here

endmodule
