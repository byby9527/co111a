`ifndef not_nt
   `include "not_nt.v"
`endif
`define or_nt 1

module or_nt(input a, input b, output out);

    // Put your code here

endmodule
