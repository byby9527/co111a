`ifndef not_nt
   `include "not_nt.v"
`endif
`define not_16 1

module not_16(
    input [15:0] in,
    output [15:0] out
);

    // Put your code here

endmodule
