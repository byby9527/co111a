`ifndef or_nt
  `include "or_nt.v"
`endif
`define or8way 1

module or8way(
    input [7:0] in,
    output      out
);

    // Put your code here

endmodule
