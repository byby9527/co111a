`ifndef half_adder
  `include "half_adder.v"
`endif
`define inc_16 1

module inc_16(input [15:0] in, output [15:0] out);

    // Put your code here  

endmodule
