`ifndef full_adder
   `include "full_adder.v"
`endif
`define add_16 1

module add_16(
    input  [15:0] a,
    input  [15:0] b,
    output [15:0] out
);

    // Put your code here
    
endmodule
