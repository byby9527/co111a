`define not_nt 1

module not_nt(input in, output out);
    
    // Put your code here

endmodule
