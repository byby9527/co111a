`ifndef and_nt
  `include "and_nt.v"
`endif
`define mux 1

module mux(
    input  a,
    input  b,
    input  select,
    output out
);

    // Put your code here

endmodule
