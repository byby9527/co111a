`ifndef or_n2t
  `include "or_n2t.sv"
`endif
`define or_8_way 1

module or_8_way(
    input [7:0] in,
    output      out
);

    // Put your code here

endmodule
