`ifndef xor_nt
  `include "../01/xor_nt.v"
`endif
`define half_adder 1

module half_adder(
    input  a,
    input  b,
    output carry,
    output sum
);

    // Put your code here

endmodule
