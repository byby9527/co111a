`ifndef and_nt
  `include "and_nt.v"
`endif
`define xor_nt 1

module xor_nt(input a, input b, output out);

    // Put your code here

endmodule
