`ifndef or_nt
  `include "or_nt.v"
`endif
`define or_16 1

module or_16(
    input[15:0] a,
    input[15:0] b,
    output[15:0] out
);

    // Put your code here

endmodule
