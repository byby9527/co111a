`ifndef or_nt
  `include "or_nt.v"
`endif
`define and_n2t 1

module and_n2t(input a, input b, output out);

    // Put your code here

endmodule 
