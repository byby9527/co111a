`ifndef and_nt
  `include "and_nt.sv"
`endif
`define dmux 1

module dmux(
    input  in,
    input  select,
    output a,
    output b
);

    // Put your code here

endmodule
